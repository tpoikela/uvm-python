//---------------------------------------------------------------------------
// File: module_top.sv
// Created on 2020-01-08
// Tuomas Poikela, tuomas.poikela@cern.ch
//
// Description: 
//---------------------------------------------------------------------------

`timescale 1ns/1ps

module module_top(input clk, input rst);

endmodule: module_top

